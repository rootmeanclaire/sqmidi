module which_note #(
	parameter F_CLK = 12_000_000;
) (
	input wire clk,
	input wire reset,
	input audio,
	// 7-bit MIDI note value
	output reg[6:0] midi,
	// High if a note is currently being played, low otherwise
	output reg note_on
);
	// Magic numbers generated along with note period LUT
	localparam P_MAX = 'h5996;
	localparam MSB = 20;
	localparam LSB = 6;
	// Timer for the current 
	reg[20:0] period = 0;

	always @(posedge reset) begin
		period <= 0;
	end

	always @(posedge audio) begin
		if (note_on) begin
			// Lookup table for note periods
			// Generated by gen-note-lut.py
			case (period[MSB:LSB])
				15: midi <= 127;
				16: midi <= 126;
				17: midi <= 125;
				18: midi <= 124;
				19: midi <= 123;
				20: midi <= 122;
				21: midi <= 121;
				22: midi <= 120;
				24: midi <= 119;
				25: midi <= 118;
				27: midi <= 117;
				28: midi <= 116;
				30: midi <= 115;
				32: midi <= 114;
				34: midi <= 113;
				36: midi <= 112;
				38: midi <= 111;
				40: midi <= 110;
				42: midi <= 109;
				45: midi <= 108;
				47: midi <= 107;
				50: midi <= 106;
				53: midi <= 105;
				56: midi <= 104;
				60: midi <= 103;
				63: midi <= 102;
				67: midi <= 101;
				71: midi <= 100;
				75: midi <= 99;
				80: midi <= 98;
				85: midi <= 97;
				90: midi <= 96;
				95: midi <= 95;
				101: midi <= 94;
				107: midi <= 93;
				113: midi <= 92;
				120: midi <= 91;
				127: midi <= 90;
				134: midi <= 89;
				142: midi <= 88;
				151: midi <= 87;
				160: midi <= 86;
				169: midi <= 85;
				179: midi <= 84;
				190: midi <= 83;
				201: midi <= 82;
				213: midi <= 81;
				226: midi <= 80;
				239: midi <= 79;
				253: midi <= 78;
				268: midi <= 77;
				284: midi <= 76;
				301: midi <= 75;
				319: midi <= 74;
				338: midi <= 73;
				358: midi <= 72;
				380: midi <= 71;
				402: midi <= 70;
				426: midi <= 69;
				451: midi <= 68;
				478: midi <= 67;
				507: midi <= 66;
				537: midi <= 65;
				569: midi <= 64;
				603: midi <= 63;
				638: midi <= 62;
				676: midi <= 61;
				717: midi <= 60;
				759: midi <= 59;
				804: midi <= 58;
				852: midi <= 57;
				903: midi <= 56;
				957: midi <= 55;
				1014: midi <= 54;
				1074: midi <= 53;
				1138: midi <= 52;
				1205: midi <= 51;
				1277: midi <= 50;
				1353: midi <= 49;
				1433: midi <= 48;
				1519: midi <= 47;
				1609: midi <= 46;
				1705: midi <= 45;
				1806: midi <= 44;
				1913: midi <= 43;
				2027: midi <= 42;
				2148: midi <= 41;
				2275: midi <= 40;
				2411: midi <= 39;
				2554: midi <= 38;
				2706: midi <= 37;
				2867: midi <= 36;
				3037: midi <= 35;
				3218: midi <= 34;
				3409: midi <= 33;
				3612: midi <= 32;
				3827: midi <= 31;
				4054: midi <= 30;
				4295: midi <= 29;
				4551: midi <= 28;
				4821: midi <= 27;
				5108: midi <= 26;
				5412: midi <= 25;
				5733: midi <= 24;
				6074: midi <= 23;
				6436: midi <= 22;
				6818: midi <= 21;
				7224: midi <= 20;
				7653: midi <= 19;
				8108: midi <= 18;
				8590: midi <= 17;
				9101: midi <= 16;
				9642: midi <= 15;
				10216: midi <= 14;
				10823: midi <= 13;
				11467: midi <= 12;
				12149: midi <= 11;
				12871: midi <= 10;
				13636: midi <= 9;
				14447: midi <= 8;
				15306: midi <= 7;
				16216: midi <= 6;
				17181: midi <= 5;
				18202: midi <= 4;
				19285: midi <= 3;
				20431: midi <= 2;
				21646: midi <= 1;
				22934: midi <= 0;
				default: note_on <= 1'b0;
			endcase
		end else begin
			note_on <= 1'b1;
		end
		period <= 0;
	end
	always @(posedge clk) begin
		period += 1;
	end
endmodule
